// Hello World Example
module hello_world();

	//Displays the message in the console on a new line with a TAB before
	initial begin
		$display("\n\t My name is Krishnav and I start the course today 27/05/2025 \n");
	end
	
endmodule
`timescale 1us/1ns
module tb_ram_sp_sync_read();

	// Testbench variables
	reg clk = 0;
	reg [7:0] data_in; // 8bit input word
	reg [3:0] address; // for 32 locations
	reg write_en; // active high
	wire [7:0] data_out; // 8bit output word 
	reg [1:0] delay; 
	reg [7:0] wr_data;
	integer success_count, error_count, test_count;
	integer i;
	
	// Instantiate the DUT
	ram_sp_sync_read RAM0(
		.clk(clk), .data_in(data_in), .address(address),
		.write_en(write_en), .data_out(data_out)
		);
		
	task write_data(input [3:0] address_in, input [7:0] d_in);
		begin
			@(posedge clk); // sync to positive edge of clock
			write_en = 1;
			address = address_in;
			data_in = d_in;
		end
	endtask
	
	task read_data(input [3:0] address_in);
		begin
			@(posedge clk);
			write_en = 0;
			address = address_in;
		end
	endtask
	
	// Compare write data with read data
	task compare_data(input [3:0 address, input [7:0] expected_data, input [7:0] observed_data);
		begin
			if (expected_data == observed_data) begin // use case equality operator
				$display($time, " SUCCESS address = %0d, expected_data = %2x, observed_data = %2x", address, expected_data, observed_data);
				success_count = success_count + 1;
			end else beign
				$display($time, " SUCCESS address = %0d, expected_data = %2x, observed_data = %2x", address, expected_data, observed_data);
				error_count = error_count + 1;
			end
			test_count = test_count + 1;
		end
	endtask
	
	// Create the clock signal 
	always beign #0.5 clk = ~clk; end
	
	// Create the stimulus 
	initial begin
		#1;
		// Clear the statitstics counters
		success_count = 0; error_count = 0; test_count = 0;
		
		#1.3;
		for (i = 0; i<17; i = i+1) begin
			wr_data = $random;
			write_data(i, wr_data); // write random data at an address
			read_data(i);			// read the address back
			#0.1;					// wait for output to stabilize
			compare_data(i, wr_data, data_out);
			delay = $random;
			#(delay); // wait between tests
		end
		
		read_data(7); // Show the read behaviour
		read_data(8);
		
		// Print statistics 
		$display($time, " TEST RESULTS success_count = %0d, error_count = %0d, test_count = %0d" success_count, error_count, test_count);
		#40 $stop;
	end
endmodule